`ifndef GON_APB_DEFINES_SVH
`define GON_APB_DEFINES_SVH

`define APB_ADDR_WIDTH 32

`endif
