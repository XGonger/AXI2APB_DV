`ifndef GON_AXI2APB_TESTS_SVH
`define GON_AXI2APB_TESTS_SVH

`include "gon_axi2apb_base_test.sv"
`include "gon_axi2apb_smoke_test.sv"

`endif
