`ifndef GON_AXI2APB_ELEM_SEQS_SVH
`define GON_AXI2APB_ELEM_SEQS_SVH

`include "gon_axi2apb_base_elem_seq.sv"
`include "gon_axi2apb_clk_reset_set_seq.sv"
`include "gon_axi2apb_write_seq.sv"
`include "gon_axi2apb_read_seq.sv"

`endif 
