`ifndef GON_AXI_SEQ_LIB_SV
`define GON_AXI_SEQ_LIB_SV

`include "gon_axi_base_seq.sv"
`include "gon_axi_transfer_seq.sv"

`endif
