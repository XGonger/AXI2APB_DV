`ifndef GON_CLK_RESET_IF_SV
`define GON_CLK_RESET_IF_SV

interface gon_clk_reset_if;
  logic clk;
  logic reset_;

endinterface


`endif
