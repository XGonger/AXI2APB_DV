`ifndef GON_APB_PKG_SV
`define GON_APB_PKG_SV

package gon_apb_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "gon_apb_defines.svh"
  `include "gon_apb_types.sv"
  `include "gon_apb_agent_configuration.sv"
  `include "gon_apb_transaction.sv"  
  `include "gon_apb_sequencer.sv"  
  `include "gon_apb_driver.sv"  
  `include "gon_apb_monitor.sv"  
  `include "gon_apb_slave_driver.sv"  
  `include "gon_apb_slave_monitor.sv"  
  `include "gon_apb_slave_sequencer.sv"  
  `include "gon_apb_slave_agent.sv"  
  `include "./sequence_lib/gon_apb_sequence_lib.svh"  

endpackage


`endif // GON_APB_PKG_SV
