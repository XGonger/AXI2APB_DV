`ifndef GON_APB_SEQUENCE_LIB_SVH
`define GON_APB_SEQUENCE_LIB_SVH

`include "gon_apb_base_sequence.sv"
`include "gon_apb_slave_ready.sv"

`endif // GON_APB_SEQUENCE_LIB_SVH
