`ifndef GON_AXI2APB_SEQ_LIB_SVH
`define GON_AXI2APB_SEQ_LIB_SVH

`include "gon_axi2apb_elem_seqs.svh"
`include "gon_axi2apb_base_virt_seq.sv"
`include "gon_axi2apb_smoke_virt_seq.sv"
`include "gon_axi2apb_free_reset_state_check_virt_seq.sv"
`include "gon_axi2apb_busy_reset_state_check_virt_seq.sv"

`endif
